module dff
